library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- btn connected to up/down pushbuttons for now but
-- eventually will get data from UART

entity game_over_display is
    port(
        clk, reset: in std_logic;
        pixel_x, pixel_y: in std_logic_vector(9 downto 0);
        life_cnt: in std_logic_vector(1 downto 0);
        graph_rgb: out std_logic_vector(2 downto 0)
    );
end game_over_display;

architecture arch of game_over_display is
    signal pix_x, pix_y: unsigned(9 downto 0);

    constant LETTER_SIZE: unsigned := to_unsigned(32, 10);
    constant LETTER_RGB: std_logic_vector := "110";

    type letter_type is array (0 to 31) of std_logic_vector(31 downto 0);

    constant G_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "11111111111111111100000000000011",
        "11111111111111111100000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111"
    );

    constant G_X_L1: unsigned := to_unsigned(220, 10);
    constant G_X_R1: unsigned := G_X_L1 + LETTER_SIZE - 1;
    constant G_Y_T1: unsigned := to_unsigned(150, 10);
    constant G_Y_B1: unsigned := G_Y_T1 + LETTER_SIZE - 1;

    signal G_rom_addr1, G_rom_col1: unsigned(4 downto 0);
    signal G_rom_data1: std_logic_vector(31 downto 0);
    signal G_rom_bit1: std_logic;

    signal sq_G_on1: std_logic;
    signal G_G_on1: std_logic;

    constant A_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011"
    );

    constant A_X_L1: unsigned := to_unsigned(260, 10);
    constant A_X_R1: unsigned := A_X_L1 + LETTER_SIZE - 1;
    constant A_Y_T1: unsigned := to_unsigned(150, 10);
    constant A_Y_B1: unsigned := A_Y_T1 + LETTER_SIZE - 1;

    signal A_rom_addr1, A_rom_col1: unsigned(4 downto 0);
    signal A_rom_data1: std_logic_vector(31 downto 0);
    signal A_rom_bit1: std_logic;

    signal sq_A_on1: std_logic;
    signal A_A_on1: std_logic;


    constant M_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011",
        "11000000000000011000000000000011"
    );

    constant M_X_L1: unsigned := to_unsigned(300, 10);
    constant M_X_R1: unsigned := M_X_L1 + LETTER_SIZE - 1;
    constant M_Y_T1: unsigned := to_unsigned(150, 10);
    constant M_Y_B1: unsigned := M_Y_T1 + LETTER_SIZE - 1;

    signal M_rom_addr1, M_rom_col1: unsigned(4 downto 0);
    signal M_rom_data1: std_logic_vector(31 downto 0);
    signal M_rom_bit1: std_logic;

    signal sq_M_on1: std_logic;
    signal M_M_on1: std_logic;


    constant E_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "00000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111"
    );

    constant E_X_L1: unsigned := to_unsigned(340, 10);
    constant E_X_R1: unsigned := E_X_L1 + LETTER_SIZE - 1;
    constant E_Y_T1: unsigned := to_unsigned(150, 10);
    constant E_Y_B1: unsigned := E_Y_T1 + LETTER_SIZE - 1;

    signal E_rom_addr1, E_rom_col1: unsigned(4 downto 0);
    signal E_rom_data1: std_logic_vector(31 downto 0);
    signal E_rom_bit1: std_logic;

    signal sq_E_on1: std_logic;
    signal E_E_on1: std_logic;

    constant E_X_L2: unsigned := to_unsigned(490, 10);
    constant E_X_R2: unsigned := E_X_L2 + LETTER_SIZE - 1;
    constant E_Y_T2: unsigned := to_unsigned(150, 10);
    constant E_Y_B2: unsigned := E_Y_T2 + LETTER_SIZE - 1;

    signal E_rom_addr2, E_rom_col2: unsigned(4 downto 0);
    signal E_rom_data2: std_logic_vector(31 downto 0);
    signal E_rom_bit2: std_logic;

    signal sq_E_on2: std_logic;
    signal E_E_on2: std_logic;


    constant O_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111"
    );

    constant O_X_L1: unsigned := to_unsigned(410, 10);
    constant O_X_R1: unsigned := O_X_L1 + LETTER_SIZE - 1;
    constant O_Y_T1: unsigned := to_unsigned(150, 10);
    constant O_Y_B1: unsigned := O_Y_T1 + LETTER_SIZE - 1;

    signal O_rom_addr1, O_rom_col1: unsigned(4 downto 0);
    signal O_rom_data1: std_logic_vector(31 downto 0);
    signal O_rom_bit1: std_logic;

    signal sq_O_on1: std_logic;
    signal O_O_on1: std_logic;


    constant V_ROM: letter_type:= (
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "01100000000000000000000000000011",
        "01100000000000000000000000000011",
        "00110000000000000000000000000110",
        "00110000000000000000000000000110",
        "00011000000000000000000000001100",
        "00011000000000000000000000001100",
        "00001100000000000000000000011000",
        "00001100000000000000000000011000",
        "00000110000000000000000000110000",
        "00000110000000000000000000110000",
        "00000011000000000000000001100000",
        "00000011000000000000000001100000",
        "00000001100000000000000011000000",
        "00000001100000000000000011000000",
        "00000000110000000000000110000000",
        "00000000110000000000000110000000",
        "00000000011000000000001100000000",
        "00000000011000000000001100000000",
        "00000000001100000000011000000000",
        "00000000001100000000011000000000",
        "00000000000110000000110000000000",
        "00000000000110000000110000000000",
        "00000000000011000001100000000000",
        "00000000000011000001100000000000",
        "00000000000001100011000000000000",
        "00000000000001100011000000000000",
        "00000000000000110110000000000000",
        "00000000000000110110000000000000",
        "00000000000000111100000000000000",
        "00000000000000111100000000000000"
    );

    constant V_X_L1: unsigned := to_unsigned(450, 10);
    constant V_X_R1: unsigned := V_X_L1 + LETTER_SIZE - 1;
    constant V_Y_T1: unsigned := to_unsigned(150, 10);
    constant V_Y_B1: unsigned := V_Y_T1 + LETTER_SIZE - 1;

    signal V_rom_addr1, V_rom_col1: unsigned(4 downto 0);
    signal V_rom_data1: std_logic_vector(31 downto 0);
    signal V_rom_bit1: std_logic;

    signal sq_V_on1: std_logic;
    signal V_V_on1: std_logic;


    constant R_ROM: letter_type:= (
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11000000000000000000000000000011",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "11111111111111111111111111111111",
        "00000000000000000000000000011011",
        "00000000000000000000000001110011",
        "00000000000000000000000111000011",
        "00000000000000000000011100000011",
        "00000000000000000001110000000011",
        "00000000000000000111000000000011",
        "00000000000000011100000000000011",
        "00000000000001110000000000000011",
        "00000000000111000000000000000011",
        "00000000011100000000000000000011",
        "00000001110000000000000000000011",
        "00000111000000000000000000000011",
        "00011100000000000000000000000011",
        "01110000000000000000000000000011",
        "11100000000000000000000000000011",
        "11100000000000000000000000000011"
    );

    constant R_X_L1: unsigned := to_unsigned(530, 10);
    constant R_X_R1: unsigned := R_X_L1 + LETTER_SIZE - 1;
    constant R_Y_T1: unsigned := to_unsigned(150, 10);
    constant R_Y_B1: unsigned := R_Y_T1 + LETTER_SIZE - 1;

    signal R_rom_addr1, R_rom_col1: unsigned(4 downto 0);
    signal R_rom_data1: std_logic_vector(31 downto 0);
    signal R_rom_bit1: std_logic;

    signal sq_R_on1: std_logic;
    signal R_R_on1: std_logic;
    
begin
    pix_x <= unsigned(pixel_x);
    pix_y <= unsigned(pixel_y);

    sq_G_on1 <= '1' when (G_X_L1 <= pix_x) and (pix_x <= G_X_R1) and (G_Y_T1 <= pix_y) and (pix_y <= G_Y_B1) else '0';
    G_rom_addr1 <= pix_y(4 downto 0) - G_Y_T1(4 downto 0);
    G_rom_col1 <= pix_x(4 downto 0) - G_X_L1(4 downto 0);
    G_rom_data1 <= G_ROM(to_integer(G_rom_addr1));
    G_rom_bit1 <= G_rom_data1(to_integer(G_rom_col1));
    G_G_on1 <= '1' when (sq_G_on1 = '1') and (G_rom_bit1 = '1') else '0';

    sq_A_on1 <= '1' when (A_X_L1 <= pix_x) and (pix_x <= A_X_R1) and (A_Y_T1 <= pix_y) and (pix_y <= A_Y_B1) else '0';
    A_rom_addr1 <= pix_y(4 downto 0) - A_Y_T1(4 downto 0);
    A_rom_col1 <= pix_x(4 downto 0) - A_X_L1(4 downto 0);
    A_rom_data1 <= A_ROM(to_integer(A_rom_addr1));
    A_rom_bit1 <= A_rom_data1(to_integer(A_rom_col1));
    A_A_on1 <= '1' when (sq_A_on1 = '1') and (A_rom_bit1 = '1') else '0';

    sq_M_on1 <= '1' when (M_X_L1 <= pix_x) and (pix_x <= M_X_R1) and (M_Y_T1 <= pix_y) and (pix_y <= M_Y_B1) else '0';
    M_rom_addr1 <= pix_y(4 downto 0) - M_Y_T1(4 downto 0);
    M_rom_col1 <= pix_x(4 downto 0) - M_X_L1(4 downto 0);
    M_rom_data1 <= M_ROM(to_integer(M_rom_addr1));
    M_rom_bit1 <= M_rom_data1(to_integer(M_rom_col1));
    M_M_on1 <= '1' when (sq_M_on1 = '1') and (M_rom_bit1 = '1') else '0';

    sq_E_on1 <= '1' when (E_X_L1 <= pix_x) and (pix_x <= E_X_R1) and (E_Y_T1 <= pix_y) and (pix_y <= E_Y_B1) else '0';
    E_rom_addr1 <= pix_y(4 downto 0) - E_Y_T1(4 downto 0);
    E_rom_col1 <= pix_x(4 downto 0) - E_X_L1(4 downto 0);
    E_rom_data1 <= E_ROM(to_integer(E_rom_addr1));
    E_rom_bit1 <= E_rom_data1(to_integer(E_rom_col1));
    E_E_on1 <= '1' when (sq_E_on1 = '1') and (E_rom_bit1 = '1') else '0';

    sq_O_on1 <= '1' when (O_X_L1 <= pix_x) and (pix_x <= O_X_R1) and (O_Y_T1 <= pix_y) and (pix_y <= O_Y_B1) else '0';
    O_rom_addr1 <= pix_y(4 downto 0) - O_Y_T1(4 downto 0);
    O_rom_col1 <= pix_x(4 downto 0) - O_X_L1(4 downto 0);
    O_rom_data1 <= O_ROM(to_integer(O_rom_addr1));
    O_rom_bit1 <= O_rom_data1(to_integer(O_rom_col1));
    O_O_on1 <= '1' when (sq_O_on1 = '1') and (O_rom_bit1 = '1') else '0';

    sq_V_on1 <= '1' when (V_X_L1 <= pix_x) and (pix_x <= V_X_R1) and (V_Y_T1 <= pix_y) and (pix_y <= V_Y_B1) else '0';
    V_rom_addr1 <= pix_y(4 downto 0) - V_Y_T1(4 downto 0);
    V_rom_col1 <= pix_x(4 downto 0) - V_X_L1(4 downto 0);
    V_rom_data1 <= V_ROM(to_integer(V_rom_addr1));
    V_rom_bit1 <= V_rom_data1(to_integer(V_rom_col1));
    V_V_on1 <= '1' when (sq_V_on1 = '1') and (V_rom_bit1 = '1') else '0';

    sq_E_on2 <= '1' when (E_X_L2 <= pix_x) and (pix_x <= E_X_R2) and (E_Y_T2 <= pix_y) and (pix_y <= E_Y_B2) else '0';
    E_rom_addr2 <= pix_y(4 downto 0) - E_Y_T2(4 downto 0);
    E_rom_col2 <= pix_x(4 downto 0) - E_X_L2(4 downto 0);
    E_rom_data2 <= E_ROM(to_integer(E_rom_addr2));
    E_rom_bit2 <= E_rom_data1(to_integer(E_rom_col2));
    E_E_on2 <= '1' when (sq_E_on2 = '1') and (E_rom_bit2 = '1') else '0';

    sq_R_on1 <= '1' when (R_X_L1 <= pix_x) and (pix_x <= R_X_R1) and (R_Y_T1 <= pix_y) and (pix_y <= R_Y_B1) else '0';
    R_rom_addr1 <= pix_y(4 downto 0) - R_Y_T1(4 downto 0);
    R_rom_col1 <= pix_x(4 downto 0) - R_X_L1(4 downto 0);
    R_rom_data1 <= R_ROM(to_integer(R_rom_addr1));
    R_rom_bit1 <= R_rom_data1(to_integer(R_rom_col1));
    R_R_on1 <= '1' when (sq_R_on1 = '1') and (R_rom_bit1 = '1') else '0';

    graph_rgb <= LETTER_RGB when ((G_G_on1 = '1') or (A_A_on1 = '1') or (M_M_on1 = '1') or (E_E_on1 = '1') or (O_O_on1 = '1') or (V_V_on1 = '1') or (E_E_on2 = '1') or (R_R_on1 = '1')) else "000";
end arch;














